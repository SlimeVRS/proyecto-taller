module n_not (output logic c, input logic a);
not operator(c,a);
endmodule