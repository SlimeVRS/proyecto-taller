module or_mux (output logic out,input logic op0000,op0001,op0010,op0011,op0100,op0101,op1000,op1001,op1010,op1011,op1100,op1101);
	or out_mux(out,op0000,op0001,op0010,op0011,op0100,op0101,op1000,op1001,op1010,op1011,op1100,op1101);
endmodule