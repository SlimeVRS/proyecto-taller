module n_xor (output logic c, input logic a,b);
	xor
		operator(c,a,b);
endmodule