module n_or (output logic C,input logic A,B);
	or operator(C,A,B);
endmodule
