module n_and(output logic c,input logic a,b);
and operator(c,a,b);
endmodule